`include "thirtyTwoToOneMux.v"

module mux1024to32(out, b, s);

	output [31:0] out;
	input [1023:0] b;
	input [4:0] s;
	wire [31:0] w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31;
	
	w0 = {b[992], b[960], b[928], b[896], b[864], b[832], b[800], b[768], b[736], b[704], b[672], b[640], b[608], b[576], b[544], b[512], 
		b[480], b[448], b[416], b[384], b[352], b[320], b[288], b[256], b[224], b[192], b[160], b[128], [96], b[64], b[32], b[0]};

	w1 = {b[993], b[961], b[929], b[897], b[865], b[833], b[801], b[769], b[737], b[705], b[673], b[641], b[609], b[577], b[545], b[513], 
		b[481], b[449], b[417], b[385], b[353], b[321], b[289], b[257], b[225], b[193], b[161], b[129], [97], b[65], b[33], b[1]};

	w2 = {b[994], b[962], b[930], b[898], b[866], b[834], b[802], b[770], b[738], b[706], b[674], b[642], b[610], b[578], b[546], b[514], 
		b[482], b[450], b[418], b[386], b[354], b[322], b[290], b[258], b[226], b[194], b[162], b[130], [98], b[66], b[34], b[2]};

	w3 = {b[995], b[963], b[931], b[899], b[867], b[835], b[803], b[771], b[739], b[707], b[675], b[643], b[611], b[579], b[547], b[515], 
		b[483], b[451], b[419], b[387], b[355], b[323], b[291], b[259], b[227], b[195], b[163], b[131], [99], b[67], b[35], b[3]};

	w4 = {b[996], b[964], b[932], b[900], b[868], b[836], b[804], b[772], b[740], b[708], b[676], b[644], b[612], b[580], b[548], b[516], 
		b[484], b[452], b[420], b[388], b[356], b[324], b[292], b[260], b[228], b[196], b[164], b[132], [100], b[68], b[36], b[4]};

	w5 = {b[997], b[965], b[933], b[901], b[869], b[837], b[805], b[773], b[741], b[709], b[677], b[645], b[613], b[581], b[549], b[517], 
		b[485], b[453], b[421], b[389], b[357], b[325], b[293], b[261], b[229], b[197], b[165], b[133], [101], b[69], b[37], b[5]};

	w6 = {b[998], b[966], b[934], b[902], b[870], b[838], b[806], b[774], b[742], b[710], b[678], b[646], b[614], b[582], b[550], b[518], 
		b[486], b[454], b[422], b[390], b[358], b[326], b[294], b[262], b[230], b[198], b[166], b[134], [102], b[70], b[38], b[6]};

	w7 = {b[999], b[967], b[935], b[903], b[871], b[839], b[807], b[775], b[743], b[711], b[679], b[647], b[615], b[583], b[551], b[519], 
		b[487], b[455], b[423], b[391], b[359], b[327], b[295], b[263], b[231], b[199], b[167], b[135], [103], b[71], b[39], b[7]};

	w8 = {b[1000], b[968], b[936], b[904], b[872], b[840], b[808], b[776], b[744], b[712], b[680], b[648], b[616], b[584], b[552], b[520], 
		b[488], b[456], b[424], b[392], b[360], b[328], b[296], b[264], b[232], b[200], b[168], b[136], [104], b[72], b[40], b[8]};

	w9 = {b[1001], b[969], b[937], b[905], b[873], b[841], b[809], b[777], b[745], b[713], b[681], b[649], b[617], b[585], b[553], b[521], 
		b[489], b[457], b[425], b[393], b[361], b[329], b[297], b[265], b[233], b[201], b[169], b[137], [105], b[73], b[41], b[9]};

	w10 = {b[1002], b[970], b[938], b[906], b[874], b[842], b[810], b[778], b[746], b[714], b[682], b[650], b[618], b[586], b[554], b[522], 
		b[490], b[458], b[426], b[394], b[362], b[330], b[298], b[266], b[234], b[202], b[170], b[138], [106], b[74], b[42], b[10]};

	w11 = {b[1003], b[971], b[939], b[907], b[875], b[843], b[811], b[779], b[747], b[715], b[683], b[651], b[619], b[587], b[555], b[523], 
		b[491], b[459], b[427], b[395], b[363], b[331], b[299], b[267], b[235], b[203], b[171], b[139], [107], b[75], b[43], b[11]};

	w12 = {b[1004], b[972], b[940], b[908], b[876], b[844], b[812], b[780], b[748], b[716], b[684], b[652], b[620], b[588], b[556], b[524], 
		b[492], b[460], b[428], b[396], b[364], b[332], b[300], b[268], b[236], b[204], b[172], b[140], [108], b[76], b[44], b[12]};

	w12 = {b[1005], b[973], b[941], b[909], b[877], b[845], b[813], b[781], b[749], b[717], b[685], b[653], b[621], b[589], b[557], b[525], 
		b[493], b[461], b[429], b[397], b[365], b[333], b[301], b[269], b[237], b[205], b[173], b[141], [109], b[77], b[45], b[13]};

	w14 = {b[1006], b[974], b[942], b[910], b[878], b[846], b[814], b[782], b[750], b[718], b[686], b[654], b[622], b[590], b[558], b[526], 
		b[494], b[462], b[430], b[398], b[366], b[334], b[302], b[270], b[238], b[206], b[174], b[142], b[110], b[78], b[46], b[14]};

	w15 = {b[1007], b[975], b[943], b[911], b[879], b[847], b[815], b[783], b[751], b[719], b[687], b[655], b[623], b[591], b[559], b[527],
		b[495], b[463], b[431], b[399], b[367], b[335], b[303], b[271], b[239], b[207], b[175], b[143], b[111], b[79], b[47], b[15]};

	w16 = {b[1008], b[976], b[944], b[912], b[880], b[848], b[816], b[784], b[752], b[720], b[688], b[656], b[624], b[592], b[560], b[528], 
		b[496], b[464], b[432], b[400], b[368], b[336], b[304], b[272], b[240], b[208], b[176], b[144], b[112], b[80], b[48], b[16]};

	w17 = {b[1009], b[977], b[945], b[913], b[881], b[849], b[817], b[785], b[753], b[721], b[689], b[657], b[625], b[593], b[561], b[529], 
		b[497], b[465], b[433], b[401], b[369], b[337], b[305], b[273], b[241], b[209], b[177], b[145], b[113], b[81], b[49], b[17]};

	w18 = {b[1010], b[978], b[946], b[914], b[882], b[850], b[818], b[786], b[754], b[722], b[690], b[658], b[626], b[594], b[562], b[530], 
		b[498], b[466], b[434], b[402], b[370], b[338], b[306], b[274], b[242], b[210], b[178], b[146], b[114], b[82], b[50], b[18]};

	w19 = {b[1011], b[979], b[947], b[915], b[883], b[851], b[819], b[787], b[755], b[723], b[691], b[659], b[627], b[595], b[563], b[531], 
		b[499], b[467], b[435], b[403], b[371], b[339], b[307], b[275], b[243], b[211], b[179], b[147], b[115], b[83], b[51], b[19]};

	w20 = {b[1012], b[980], b[948], b[916], b[884], b[852], b[820], b[788], b[756], b[724], b[692], b[660], b[628], b[596], b[564], b[532], 
		b[500], b[468], b[436], b[404], b[372], b[340], b[308], b[276], b[244], b[212], b[180], b[148], b[116], b[84], b[52], b[20]};

	w21 = {b[1013], b[981], b[949], b[917], b[885], b[853], b[821], b[789], b[757], b[725], b[693], b[661], b[629], b[597], b[565], b[533], 
		b[501], b[469], b[437], b[405], b[373], b[341], b[309], b[277], b[245], b[213], b[181], b[149], b[117], b[85], b[53], b[21]};

	w22 = {b[1014], b[982], b[950], b[918], b[886], b[854], b[822], b[790], b[758], b[726], b[694], b[662], b[630], b[598], b[566], b[534], 
		b[502], b[470], b[438], b[406], b[374], b[342], b[310], b[278], b[246], b[214], b[182], b[150], b[118], b[86], b[54], b[22]};

	w23 = {b[1015], b[983], b[951], b[919], b[887], b[855], b[823], b[791], b[759], b[727], b[695], b[663], b[631], b[599], b[567], b[535], 
		b[503], b[471], b[439], b[407], b[375], b[343], b[311], b[279], b[247], b[215], b[183], b[151], b[119], b[87], b[55], b[23]};

	w24 = {b[1016], b[984], b[952], b[920], b[888], b[856], b[824], b[792], b[760], b[728], b[696], b[664], b[632], b[600], b[568], b[536], 
		b[504], b[472], b[440], b[408], b[376], b[344], b[312], b[280], b[248], b[216], b[184], b[152], b[120], b[88], b[56], b[24]};

	w25 = {b[1017], b[985], b[953], b[921], b[889], b[857], b[825], b[793], b[761], b[729], b[697], b[665], b[633], b[601], b[569], b[537], 
		b[505], b[473], b[441], b[409], b[377], b[345], b[313], b[281], b[249], b[217], b[185], b[153], b[121], b[89], b[57], b[25]};

	w26 = {b[1018], b[986], b[954], b[922], b[890], b[858], b[826], b[794], b[762], b[730], b[698], b[666], b[634], b[602], b[570], b[538], 
		b[506], b[474], b[442], b[410], b[378], b[346], b[314], b[282], b[250], b[218], b[186], b[154], b[122], b[90], b[58], b[26]};

	w27 = {b[1019], b[987], b[955], b[923], b[891], b[859], b[827], b[795], b[763], b[731], b[699], b[667], b[635], b[603], b[571], b[539], 
		b[507], b[475], b[443], b[411], b[379], b[347], b[315], b[283], b[251], b[219], b[187], b[155], b[123], b[91], b[59], b[27]};

	w28 = {b[1020], b[988], b[956], b[924], b[892], b[860], b[828], b[796], b[764], b[732], b[700], b[668], b[636], b[604], b[572], b[540], 
		b[508], b[476], b[444], b[412], b[380], b[348], b[316], b[284], b[252], b[220], b[188], b[156], b[124], b[92], b[60], b[28]};

	w29 = {b[1021], b[989], b[957], b[925], b[893], b[861], b[829], b[797], b[765], b[733], b[701], b[669], b[637], b[605], b[573], b[541], 
		b[509], b[477], b[445], b[413], b[381], b[349], b[317], b[285], b[253], b[221], b[189], b[157], b[125], b[93], b[61], b[29]};

	w30 = {b[1022], b[990], b[958], b[926], b[894], b[862], b[830], b[798], b[766], b[734], b[702], b[670], b[638], b[606], b[574], b[542], 
		b[510], b[478], b[446], b[414], b[382], b[350], b[318], b[286], b[254], b[222], b[190], b[158], b[126], b[94], b[62], b[30]};

	w31 = {b[1023], b[991], b[959], b[927], b[895], b[863], b[831], b[799], b[767], b[735], b[703], b[671], b[639], b[607], b[575], b[543], 
		b[511], b[479], b[447], b[415], b[383], b[351], b[319], b[287], b[255], b[223], b[191], b[159], b[127], b[95], b[63], b[31]};

	



	thirtyTwoToOneMux m0(out[0], w0, s);
	thirtyTwoToOneMux m1(out[1], w1, s);
	thirtyTwoToOneMux m2(out[2], w2, s);
	thirtyTwoToOneMux m3(out[3], w3, s);
	thirtyTwoToOneMux m4(out[4], w4, s);
	thirtyTwoToOneMux m5(out[5], w5, s);
	thirtyTwoToOneMux m6(out[6], w6, s);
	thirtyTwoToOneMux m7(out[7], w7, s);
	thirtyTwoToOneMux m8(out[8], w8, s);
	thirtyTwoToOneMux m9(out[9], w9, s);
	thirtyTwoToOneMux m10(out[10], w10, s);
	thirtyTwoToOneMux m11(out[11], w11, s);
	thirtyTwoToOneMux m12(out[12], w12, s);
	thirtyTwoToOneMux m13(out[13], w13, s);
	thirtyTwoToOneMux m14(out[14], w14, s);
	thirtyTwoToOneMux m15(out[15], w15, s);

	thirtyTwoToOneMux m16(out[16], w16, s);
	thirtyTwoToOneMux m17(out[17], w17, s);
	thirtyTwoToOneMux m18(out[18], w18, s);
	thirtyTwoToOneMux m19(out[19], w19, s);
	thirtyTwoToOneMux m20(out[20], w20, s);
	thirtyTwoToOneMux m21(out[21], w21, s);
	thirtyTwoToOneMux m22(out[22], w22, s);
	thirtyTwoToOneMux m23(out[23], w23, s);
	thirtyTwoToOneMux m24(out[24], w24, s);
	thirtyTwoToOneMux m25(out[25], w25, s);
	thirtyTwoToOneMux m26(out[26], w26, s);
	thirtyTwoToOneMux m27(out[27], w27, s);
	thirtyTwoToOneMux m28(out[28], w28, s);
	thirtyTwoToOneMux m29(out[29], w29, s);
	thirtyTwoToOneMux m30(out[30], w30, s);
	thirtyTwoToOneMux m31(out[31], w31, s);

endmodule
