`include "D_FF.v"
module thirtyTwoBitRegister(out, in, writeEnable, rst, clk);
	output [31:0] out;
	input [31:0] in;
	input writeEnable, rst, clk;
	wire [31:0] d;
	
	twoToOneMux ttoMux0(d[0], out[0], in[0], writeEnable);
	twoToOneMux ttoMux1(d[1], out[1], in[1], writeEnable);
	twoToOneMux ttoMux2(d[2], out[2], in[2], writeEnable);
	twoToOneMux ttoMux3(d[3], out[3], in[3], writeEnable);
	twoToOneMux ttoMux4(d[4], out[4], in[4], writeEnable);
	twoToOneMux ttoMux5(d[5], out[5], in[5], writeEnable);
	twoToOneMux ttoMux6(d[6], out[6], in[6], writeEnable);
	twoToOneMux ttoMux7(d[7], out[7], in[7], writeEnable);
	twoToOneMux ttoMux8(d[8], out[8], in[8], writeEnable);
	twoToOneMux ttoMux9(d[9], out[9], in[9], writeEnable);
	twoToOneMux ttoMux10(d[10], out[10], in[10], writeEnable);
	twoToOneMux ttoMux11(d[11], out[11], in[11], writeEnable);
	twoToOneMux ttoMux12(d[12], out[12], in[12], writeEnable);
	twoToOneMux ttoMux13(d[13], out[13], in[13], writeEnable);
	twoToOneMux ttoMux14(d[14], out[14], in[14], writeEnable);
	twoToOneMux ttoMux15(d[15], out[15], in[15], writeEnable);
	twoToOneMux ttoMux16(d[16], out[16], in[16], writeEnable);
	twoToOneMux ttoMux17(d[17], out[17], in[17], writeEnable);
	twoToOneMux ttoMux18(d[18], out[18], in[18], writeEnable);
	twoToOneMux ttoMux19(d[19], out[19], in[19], writeEnable);
	twoToOneMux ttoMux20(d[20], out[20], in[20], writeEnable);
	twoToOneMux ttoMux21(d[21], out[21], in[21], writeEnable);
	twoToOneMux ttoMux22(d[22], out[22], in[22], writeEnable);
	twoToOneMux ttoMux23(d[23], out[23], in[23], writeEnable);
	twoToOneMux ttoMux24(d[24], out[24], in[24], writeEnable);
	twoToOneMux ttoMux25(d[25], out[25], in[25], writeEnable);
	twoToOneMux ttoMux26(d[26], out[26], in[26], writeEnable);
	twoToOneMux ttoMux27(d[27], out[27], in[27], writeEnable);
	twoToOneMux ttoMux28(d[28], out[28], in[28], writeEnable);
	twoToOneMux ttoMux29(d[29], out[29], in[29], writeEnable);
	twoToOneMux ttoMux30(d[30], out[30], in[30], writeEnable);
	twoToOneMux ttoMux31(d[31], out[31], in[31], writeEnable);
	D_FF bit0(out[0], d[0], rst, clk);
 	D_FF bit1(out[1], d[1], rst, clk);
	D_FF bit2(out[2], d[2], rst, clk);
	D_FF bit3(out[3], d[3], rst, clk);
	D_FF bit4(out[4], d[4], rst, clk);
	D_FF bit5(out[5], d[5], rst, clk);
	D_FF bit6(out[6], d[6], rst, clk);
	D_FF bit7(out[7], d[7], rst, clk);
	D_FF bit8(out[8], d[8], rst, clk);
	D_FF bit9(out[9], d[9], rst, clk);
	D_FF bit10(out[10], d[10], rst, clk);
	D_FF bit11(out[11], d[11], rst, clk);
	D_FF bit12(out[12], d[12], rst, clk);
	D_FF bit13(out[13], d[13], rst, clk);
	D_FF bit14(out[14], d[14], rst, clk);
	D_FF bit15(out[15], d[15], rst, clk);
	D_FF bit16(out[16], d[16], rst, clk);
	D_FF bit17(out[17], d[17], rst, clk);
	D_FF bit18(out[18], d[18], rst, clk);
	D_FF bit19(out[19], d[19], rst, clk);
	D_FF bit20(out[20], d[20], rst, clk);
	D_FF bit21(out[21], d[21], rst, clk);
	D_FF bit22(out[22], d[22], rst, clk);
	D_FF bit23(out[23], d[23], rst, clk);
	D_FF bit24(out[24], d[24], rst, clk);
	D_FF bit25(out[25], d[25], rst, clk);
	D_FF bit26(out[26], d[26], rst, clk);
	D_FF bit27(out[27], d[27], rst, clk);
	D_FF bit28(out[28], d[28], rst, clk);
	D_FF bit29(out[29], d[29], rst, clk);
	D_FF bit30(out[30], d[30], rst, clk);
	D_FF bit31(out[31], d[31], rst, clk);
endmodule
