`include "fiveToThirtyTwoDecoder.v"


module testBenchDecoder();
initial
	begin
		$shm_open("waves.shm");
		$shm_probe("AC");
		$shm_close(0);
	end
	reg [4:0] w;
	reg en;
	wire [31:0] y;

   fiveToThirtyTwoDecoder FiveTo32Decoder(y, w, en);

   initial
	
     begin
	en = 1;
	#1000;
	w[0] = 0;
	w[1] = 0;
	w[2] = 0;
	w[3] = 0;
	w[4] = 0;
	#1000;
	w[0] = 1;
	w[1] = 0;
	w[2] = 0;
	w[3] = 0;
	w[4] = 0;
	#1000;
	w[0] = 0;
	w[1] = 1;
	w[2] = 0;
	w[3] = 0;
	w[4] = 0;

	#1000;
	w[0] = 1;
	w[1] = 1;
	w[2] = 0;
	w[3] = 0;
	w[4] = 0;
	#1000;
	w[0] = 0;
	w[1] = 0;
	w[2] = 1;
	w[3] = 0;
	w[4] = 0;
	#1000;
	w[0] = 1;
	w[1] = 0;
	w[2] = 1;
	w[3] = 0;
	w[4] = 0;
	#1000;
	w[0] = 0;
	w[1] = 1;
	w[2] = 1;
	w[3] = 0;
	w[4] = 0;
	#1000;
	w[0] = 1;
	w[1] = 1;
	w[2] = 1;
	w[3] = 0;
	w[4] = 0;
	#1000;
	w[0] = 0;
	w[1] = 0;
	w[2] = 0;
	w[3] = 1;
	w[4] = 0;
	#1000;
	w[0] = 1;
	w[1] = 0;
	w[2] = 0;
	w[3] = 1;
	w[4] = 0;
	#1000;
	w[0] = 0;
	w[1] = 1;
	w[2] = 0;
	w[3] = 1;
	w[4] = 0;
	#1000;
	w[0] = 1;
	w[1] = 1;
	w[2] = 0;
	w[3] = 1;
	w[4] = 0;
	#1000;
	w[0] = 0;
	w[1] = 0;
	w[2] = 1;
	w[3] = 1;
	w[4] = 0;
	#1000;
	w[0] = 1;
	w[1] = 0;
	w[2] = 1;
	w[3] = 1;
	w[4] = 0;
	#1000;
	w[0] = 0;
	w[1] = 1;
	w[2] = 1;
	w[3] = 1;
	w[4] = 0;
	#1000;
	w[0] = 1;
	w[1] = 1;
	w[2] = 1;
	w[3] = 1;
	w[4] = 0;
	#1000;
	w[0] = 0;
	w[1] = 1;
	w[2] = 1;
	w[3] = 1;
	w[4] = 1;
	#1000;
	w[0] = 1;
	w[1] = 1;
	w[2] = 1;
	w[3] = 1;
	w[4] = 1;
     end // initial begin
endmodule // testBenchDecoder

   
