module norFunct(out, in1, in2);
	output [31:0] out;
	input [31:0] in1, in2;

	nor a(out[0], in1[0], in2[0]);
	nor b(out[1], in1[1], in2[1]);
	nor c(out[2], in1[2], in2[2]);
	nor d(out[3], in1[3], in2[3]);
	nor e(out[4], in1[4], in2[4]);
	nor f(out[5], in1[5], in2[5]);
	nor g(out[6], in1[6], in2[6]);
	nor h(out[7], in1[7], in2[7]);
	nor i(out[8], in1[8], in2[8]);
	nor j(out[9], in1[9], in2[9]);
	nor k(out[10], in1[10], in2[10]);
	nor l(out[11], in1[11], in2[11]);
	nor m(out[12], in1[12], in2[12]);
	nor n(out[13], in1[13], in2[13]);
	nor o(out[14], in1[14], in2[14]);
	nor p(out[15], in1[15], in2[15]);
	nor q(out[16], in1[16], in2[16]);
	nor r(out[17], in1[17], in2[17]);
	nor s(out[18], in1[18], in2[18]);
	nor t(out[19], in1[19], in2[19]);
	nor u(out[20], in1[20], in2[20]);
	nor v(out[21], in1[21], in2[21]);
	nor w(out[22], in1[22], in2[22]);
	nor x(out[23], in1[23], in2[23]);
	nor y(out[24], in1[24], in2[24]);
	nor z(out[25], in1[25], in2[25]);
	nor aa(out[26], in1[26], in2[26]);
	nor ab(out[27], in1[27], in2[27]);
	nor ac(out[28], in1[28], in2[28]);
	nor ad(out[29], in1[29], in2[29]);
	nor ae(out[30], in1[30], in2[30]);
	nor af(out[31], in1[31], in2[31]);

endmodule
